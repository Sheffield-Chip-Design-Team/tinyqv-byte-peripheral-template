`default_nettype none
`timescale 1ns / 1ps

/* This testbench just instantiates the module and makes some convenient wires
   that can be driven / tested by the cocotb test.py.
*/

`ifndef VCD_PATH
  `define VCD_PATH "tb.vcd"
`endif

module tb ();

  string vcdname; 

  // Wire up the inputs and outputs:
  reg clk;
  reg rst_n;
  reg ena;
  reg [7:0] ui_in;
  reg [7:0] uio_in;
  wire [7:0] uo_out;
  wire [7:0] uio_out;
  wire [7:0] uio_oe;
`ifdef GL_TEST
  wire VPWR = 1'b1;
  wire VGND = 1'b0;
`endif

  // helper signals for testbench debug
  reg nes_latch;
  reg nes_clk;
  reg nes_data;

  always @(*) begin
    nes_latch = uo_out[6];
    nes_clk   = uo_out[7];
    ui_in[1]  = nes_data;
  end

  tt_um_tqv_peripheral_harness test_harness (

      // Include power ports for the Gate Level test:
`ifdef GL_TEST
      .VPWR(VPWR),
      .VGND(VGND),
`endif

      .ui_in  (ui_in),    // Dedicated inputs
      .uo_out (uo_out),   // Dedicated outputs
      .uio_in (uio_in),   // IOs: Input path
      .uio_out(uio_out),  // IOs: Output path
      .uio_oe (uio_oe),   // IOs: Enable path (active high: 0=input, 1=output)
      .ena    (ena),      // enable - goes high when design is selected
      .clk    (clk),      // clock
      .rst_n  (rst_n)     // not reset
  );

    initial begin
    nes_latch = 0;
    nes_clk = 0;
    nes_data = 0;
   // Dump the signals to a VCD file. You can view it with gtkwave or surfer.
    if ($value$plusargs("VCD_PATH=%s", vcdname)) begin
      $dumpfile(vcdname);
    end else begin
      $dumpfile("tb.vcd");
    end
    $dumpvars(0, tb);
    #1;
  end

endmodule
